module testCorrelation_32 # (parameter N = 32)
(
);
    reg [31:0] Num_1,Num_2,Num_3,Num_4,Num_5,Num_6,Num_7,Num_8,Num_9,Num_10,Num_11,Num_12,Num_13,Num_14,Num_15,Num_16;
    reg [31:0] Target_Num;
    reg Clock, Reset;
    wire [3:0] Out_4;
    
    Correlation_32 c(Num_1,Num_2,Num_3,Num_4,Num_5,Num_6,Num_7,Num_8,Num_9,Num_10,Num_11,Num_12,Num_13,Num_14,Num_15,Num_16,Target_Num, Clock, Reset, Out_4);

	initial begin
        Clock = 1;
        repeat(200) begin
            #5 Clock = ~Clock;
        end
    end
    initial
		begin
            $monitor("%d	\nNum_1 = %b,\nNum_2 = %b,\nNum_3 = %b,\nNum_4 = %b,\nNum_5 = %b,\nNum_6 = %b,\nNum_7 = %b,\nNum_8 = %b,\nNum_9 = %b,\nNum_10 = %b,\nNum_11 = %b,\nNum_12 = %b,\nNum_13 = %b,\nNum_14 = %b,\nNum_15 = %b,\nNum_16 = %b,\n Target_Num = %b, Clock = %b, Reset = %b, Out_4 = %b", $time,Num_1,Num_2,Num_3,Num_4,Num_5,Num_6,Num_7,Num_8,Num_9,Num_10,Num_11,Num_12,Num_13,Num_14,Num_15,Num_16, Target_Num, Clock, Reset, Out_4);
            
            Reset = 0;
            #13
            
            //Num_1 = 32'b11011011101010001110000000010011;
            Num_1 = 32'b00000000000000000000000000000000;
            Num_2 = 32'b00110110000000000101010001101010;
            Num_3 = 32'b01000110100000000110011000100111;
            Num_4 = 32'b10001111000000110000001001010111;
            Num_5 = 32'b10110010110101100100010110100000;
            Num_6 = 32'b01010101100000111111010001011011;
            Num_7 = 32'b00010001100100111100001001001000;
            Num_8 = 32'b11010011110010001100101010110001;
            Num_9 = 32'b11010100000101010011111100000001;
            Num_10 = 32'b11000010001001110110101111000110;
            Num_11 = 32'b01111010001011010010001001010111;
            Num_12 = 32'b00000100100101101100000101100010;
            Num_13 = 32'b00111101101001101110101010010111;
            Num_14 = 32'b01100111011101001110001001111101;
            Num_15 = 32'b11010011000000101010110100101000;
            Num_16 = 32'b10101011011001100111000001111110;

            Target_Num = 32'b11111111111111111111111111111111;

            #13

            //Num_1 = 32'b00010000111011101110011110101110;
            Num_1 = 32'b11111111111111111111111111111111;
            Num_2 = 32'b11001101111000000100001111010110;
            Num_3 = 32'b10010000001101111101111100001101;
            Num_4 = 32'b01010100001100101011010010111010;
            Num_5 = 32'b00101000010101111000111110111110;
            Num_6 = 32'b00100001010010110111110110110011;
            Num_7 = 32'b10110011110011001010000010111010;
            Num_8 = 32'b10001101100000100111000011101011;
            Num_9 = 32'b00010011010000110011011100111111;
            Num_10 = 32'b00011000111011000001110001010001;
            Num_11 = 32'b11110101001101100000100110100100;
            Num_12 = 32'b00010101000111110000101110001011;
            Num_13 = 32'b11101111000001101101000001000000;
            Num_14 = 32'b10111010010111010001101010111001;
            Num_15 = 32'b11000001001101001000010110011110;
            Num_16 = 32'b10101011011001100111000001111110;

            Target_Num = 32'b00000000000000000000000000000000;

            #13
            
            //Num_1 = 32'b11011011101010001110000000010011;
            Num_1 = 32'b11111111111111111111111111111111;
            Num_2 = 32'b00110110000000000101010001101010;
            Num_3 = 32'b01000110100000000110011000100111;
            Num_4 = 32'b10001111000000110000001001010111;
            Num_5 = 32'b10110010110101100100010110100000;
            Num_6 = 32'b01010101100000111111010001011011;
            Num_7 = 32'b00010001100100111100001001001000;
            Num_8 = 32'b11010011110010001100101010110001;
            Num_9 = 32'b11010100000101010011111100000001;
            Num_10 = 32'b11000010001001110110101111000110;
            Num_11 = 32'b01111010001011010010001001010111;
            Num_12 = 32'b00000100100101101100000101100010;
            Num_13 = 32'b00111101101001101110101010010111;
            Num_14 = 32'b01100111011101001110001001111101;
            Num_15 = 32'b11010011000000101010110100101000;
            Num_16 = 32'b10101011011001100111000001111110;

            Target_Num = 32'b00000000000000000000000000000000;
            
            #13

            //Num_1 = 32'b00010000111011101110011110101110;
            Num_1 = 32'b00000000000000000000000000000000;
            Num_2 = 32'b11001101111000000100001111010110;
            Num_3 = 32'b10010000001101111101111100001101;
            Num_4 = 32'b01010100001100101011010010111010;
            Num_5 = 32'b00101000010101111000111110111110;
            Num_6 = 32'b00100001010010110111110110110011;
            Num_7 = 32'b10110011110011001010000010111010;
            Num_8 = 32'b10001101100000100111000011101011;
            Num_9 = 32'b00010011010000110011011100111111;
            Num_10 = 32'b00011000111011000001110001010001;
            Num_11 = 32'b11110101001101100000100110100100;
            Num_12 = 32'b00010101000111110000101110001011;
            Num_13 = 32'b11101111000001101101000001000000;
            Num_14 = 32'b10111010010111010001101010111001;
            Num_15 = 32'b11000001001101001000010110011110;
            Num_16 = 32'b11010110011000011111100100100000;

            Target_Num = 32'b11111111111111111111111111111111;


		end
endmodule
