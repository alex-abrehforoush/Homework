
module TestSixteenThirtyTwoByOneMux;
	reg [15:0] a31, a30, a29, a28, a27, a26, a25, a24, a23, a22, a21, a20, a19, a18, a17, a16, a15, a14, a13, a12, a11, a10, a9, a8, a7, a6, a5, a4, a3, a2, a1, a0;
	reg [4:0] s;
	wire [15:0] d;
	SixteenThirtyTwoByOneMux tester(.a31(a31), .a30(a30), .a29(a29), .a28(a28), .a27(a27), .a26(a26), .a25(a25), .a24(a24), .a23(a23), .a22(a22), .a21(a21), .a20(a20), .a19(a19), .a18(a18), .a17(a17), .a16(a16), .a15(a15), .a14(a14), .a13(a13), .a12(a12), .a11(a11), .a10(a10), .a9(a9), .a8(a8), .a7(a7), .a6(a6), .a5(a5), .a4(a4), .a3(a3), .a2(a2), .a1(a1), .a0(a0), .s(s), .d(d));
	initial
		begin
			$monitor("%d	a31 = %b, a30 = %b, a29 = %b, a28 = %b, a27 = %b, a26 = %b, a25 = %b, a24 = %b, a23 = %b, a22 = %b, a21 = %b, a20 = %b, a19 = %b, a18 = %b, a17 = %b, a16 = %b, a15 = %b, a14 = %b, a13 = %b, a12 = %b, a11 = %b, a10 = %b, a9 = %b, a8 = %b, a7 = %b, a6 = %b, a5 = %b, a4 = %b, a3 = %b, a2 = %b, a1 = %b, a0 = %b, s = %b, d = %b", $time, a31, a30, a29, a28, a27, a26, a25, a24, a23, a22, a21, a20, a19, a18, a17, a16, a15, a14, a13, a12, a11, a10, a9, a8, a7, a6, a5, a4, a3, a2, a1, a0, s, d);
			
			#20
			a31 = 16'b0110001011001111;
			a30 = 16'b0101100001101100;
			a29 = 16'b0011001000000100;
			a28 = 16'b1000100010111110;
			a27 = 16'b1010100000000011;
			a26 = 16'b1101010000011101;
			a25 = 16'b1011100110101110;
			a24 = 16'b1111011001111100;
			a23 = 16'b0011100011101011;
			a22 = 16'b1101010101010001;
			a21 = 16'b1100101010110001;
			a20 = 16'b0111000110000011;
			a19 = 16'b1001110000011011;
			a18 = 16'b1011001000100111;
			a17 = 16'b1010011001000110;
			a16 = 16'b1011010001000001;
			a15 = 16'b0110110001011111;
			a14 = 16'b1001001110011000;
			a13 = 16'b0010011010001101;
			a12 = 16'b1000110110111101;
			a11 = 16'b0010000111110011;
			a10 = 16'b0100001000001101;
			a9 = 16'b0101100100010000;
			a8 = 16'b0110000010100001;
			a7 = 16'b1110111001000001;
			a6 = 16'b1101000110000111;
			a5 = 16'b1010101110011111;
			a4 = 16'b0100100111011000;
			a3 = 16'b0101101110100000;
			a2 = 16'b1100101101111000;
			a1 = 16'b1111001011010001;
			a0 = 16'b1000001000000011;
			s = 5'b01010;

			#20
			a31 = 16'b0010001011101100;
			a30 = 16'b0010000000101011;
			a29 = 16'b0011110100010111;
			a28 = 16'b1100100000101010;
			a27 = 16'b0110010011101000;
			a26 = 16'b0101111110111001;
			a25 = 16'b0000100111100111;
			a24 = 16'b1111000111000001;
			a23 = 16'b1111010001011000;
			a22 = 16'b0111101001101010;
			a21 = 16'b0001010101010101;
			a20 = 16'b0101011000001101;
			a19 = 16'b0100000010101110;
			a18 = 16'b1100110010011100;
			a17 = 16'b1010101001101000;
			a16 = 16'b0101101111000100;
			a15 = 16'b0101001011100001;
			a14 = 16'b1011101000101101;
			a13 = 16'b0111110011111000;
			a12 = 16'b0110101101011110;
			a11 = 16'b1010010001001110;
			a10 = 16'b1011001011011110;
			a9 = 16'b1100110010001111;
			a8 = 16'b1000001000011100;
			a7 = 16'b1010010011100100;
			a6 = 16'b0100011000011001;
			a5 = 16'b1000001101011111;
			a4 = 16'b1011100100111010;
			a3 = 16'b1110100101011011;
			a2 = 16'b1001010100000000;
			a1 = 16'b1100110100110011;
			a0 = 16'b0101101011100000;
			s = 5'b11001;


			#20
			a31 = 16'b0011001000000101;
			a30 = 16'b1100100101101011;
			a29 = 16'b0101101110011100;
			a28 = 16'b1011100000000110;
			a27 = 16'b1010111010001011;
			a26 = 16'b0010001111111101;
			a25 = 16'b1101010111000010;
			a24 = 16'b0110111010011101;
			a23 = 16'b0001010010100111;
			a22 = 16'b0000000011001100;
			a21 = 16'b0000100010001011;
			a20 = 16'b1011111111000110;
			a19 = 16'b0011111011111010;
			a18 = 16'b0111111101111010;
			a17 = 16'b0100011110001000;
			a16 = 16'b1100011000111110;
			a15 = 16'b1000101101101110;
			a14 = 16'b0110110100110100;
			a13 = 16'b1110011010000000;
			a12 = 16'b1111000001011111;
			a11 = 16'b0010001111100111;
			a10 = 16'b1110001001101000;
			a9 = 16'b0001010101011011;
			a8 = 16'b1011101000011100;
			a7 = 16'b0100110011111110;
			a6 = 16'b1001010011101001;
			a5 = 16'b0010101101111010;
			a4 = 16'b0010010110111100;
			a3 = 16'b0110110100100100;
			a2 = 16'b1010001000010010;
			a1 = 16'b1101010010111000;
			a0 = 16'b0000011000010101;
			s = 5'b10001;


			#20
			a31 = 16'b1100101001100110;
			a30 = 16'b1101000100011111;
			a29 = 16'b1110100001001110;
			a28 = 16'b1100101000011010;
			a27 = 16'b1110001111011010;
			a26 = 16'b1000011100010010;
			a25 = 16'b1001110110101011;
			a24 = 16'b1000010111000010;
			a23 = 16'b1100010110110000;
			a22 = 16'b1110011111001100;
			a21 = 16'b0010101101110101;
			a20 = 16'b0101001000100000;
			a19 = 16'b1110110101100000;
			a18 = 16'b0001100100111001;
			a17 = 16'b1110000110001111;
			a16 = 16'b0000101100010111;
			a15 = 16'b0000011001011111;
			a14 = 16'b0001010100000001;
			a13 = 16'b0101110110001110;
			a12 = 16'b0000001001111110;
			a11 = 16'b0011101001001000;
			a10 = 16'b0001000010010001;
			a9 = 16'b1110100001001101;
			a8 = 16'b1100011110101010;
			a7 = 16'b1110110100101111;
			a6 = 16'b0101110101111101;
			a5 = 16'b0110101000011001;
			a4 = 16'b0110110010011010;
			a3 = 16'b0011001100110000;
			a2 = 16'b1111111000111111;
			a1 = 16'b0101101001101000;
			a0 = 16'b0001101110100100;
			s = 5'b00100;
		end
endmodule